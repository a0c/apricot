library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package settings_pkg is
  type cS2_type is integer range 1 to 3;
  
end settings_pkg ;
